`timescale 1ns / 1ps

module ripplecarry4bit_stimuli(
    );
    reg [3:0]a,b;
    reg cin;
    wire [3:0]sum;
    wire cout;
    ripplecarry4bit uut(sum,cout,a,b,cin);
    initial
    begin
    a=4'b0000;b=4'b0000;cin=0;
    #10 a=4'b0000;b=4'b0000;cin=1;
    #10 a=4'b0000;b=4'b0001;cin=0;
    #10 a=4'b0000;b=4'b0001;cin=1;
    #10 a=4'b0000;b=4'b0010;cin=0;
    #10 a=4'b0000;b=4'b0010;cin=1;
    #10 a=4'b0000;b=4'b0011;cin=0;
    #10 a=4'b0000;b=4'b0011;cin=1;
    #10 a=4'b0000;b=4'b0100;cin=0;
    #10 a=4'b0000;b=4'b0100;cin=1;
    #10 a=4'b0000;b=4'b0101;cin=0;
    #10 a=4'b0000;b=4'b0101;cin=1;
    #10 a=4'b0000;b=4'b0110;cin=0;
    #10 a=4'b0000;b=4'b0110;cin=1;
    #10 a=4'b0000;b=4'b0111;cin=0;
    #10 a=4'b0000;b=4'b0111;cin=1;
    #10 a=4'b0000;b=4'b1000;cin=0;
    #10 a=4'b0000;b=4'b1000;cin=1;
    #10 a=4'b0000;b=4'b1001;cin=0;
    #10 a=4'b0000;b=4'b1001;cin=1;
    #10 a=4'b0000;b=4'b1010;cin=0;
    #10 a=4'b0000;b=4'b1010;cin=1;
    #10 a=4'b0000;b=4'b1011;cin=0;
    #10 a=4'b0000;b=4'b1011;cin=1;
    #10 a=4'b0000;b=4'b1100;cin=0;
    #10 a=4'b0000;b=4'b1100;cin=1;
    #10 a=4'b0000;b=4'b1101;cin=0;
    #10 a=4'b0000;b=4'b1101;cin=1;
    #10 a=4'b0000;b=4'b1110;cin=0;
    #10 a=4'b0000;b=4'b1110;cin=1;
    #10 a=4'b0000;b=4'b1111;cin=0;
    #10 a=4'b0000;b=4'b1111;cin=1;
 //a bits are changed from these sequence     
    #10 b=4'b1111;a=4'b0001;cin=0;
    #10 b=4'b1111;a=4'b0001;cin=1;
    #10 b=4'b1111;a=4'b0010;cin=0;
    #10 b=4'b1111;a=4'b0010;cin=1;
    #10 b=4'b1111;a=4'b0011;cin=0;
    #10 b=4'b1111;a=4'b0011;cin=1;
    #10 b=4'b1111;a=4'b0100;cin=0;
    #10 b=4'b1111;a=4'b0100;cin=1;
    #10 b=4'b1111;a=4'b0101;cin=0;
    #10 b=4'b1111;a=4'b0101;cin=1;
    #10 b=4'b1111;a=4'b0110;cin=0;
    #10 b=4'b1111;a=4'b0110;cin=1;
    #10 b=4'b1111;a=4'b0111;cin=0;
    #10 b=4'b1111;a=4'b0111;cin=1;
    #10 b=4'b1111;a=4'b1000;cin=0;
    #10 b=4'b1111;a=4'b1000;cin=1;
    #10 b=4'b1111;a=4'b1001;cin=0;
    #10 b=4'b1111;a=4'b1001;cin=1;
    #10 b=4'b1111;a=4'b1010;cin=0;
    #10 b=4'b1111;a=4'b1010;cin=1;
    #10 b=4'b1111;a=4'b1011;cin=0;
    #10 b=4'b1111;a=4'b1011;cin=1;
    #10 b=4'b1111;a=4'b1100;cin=0;
    #10 b=4'b1111;a=4'b1100;cin=1;
    #10 b=4'b1111;a=4'b1101;cin=0;
    #10 b=4'b1111;a=4'b1101;cin=1;
    #10 b=4'b1111;a=4'b1110;cin=0;
    #10 b=4'b1111;a=4'b1110;cin=1;
    #10 b=4'b1111;a=4'b1111;cin=0;
    #10 b=4'b1111;a=4'b1111;cin=1;
     
    #10 $finish;
    end    
endmodule
